library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

package song_pkg is
    type composer_song_t is (s_quiet, s_looser, s_move);

end package;
