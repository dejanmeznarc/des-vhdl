library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use work.screen_pkg.all;

entity buttons is
  port (
    clk : in std_logic
  );
end entity;
