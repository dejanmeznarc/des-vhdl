library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity control is
  port (
    clk     : in std_logic;
    buttons : in unsigned(4 downto 0)
  );
end entity;

architecture rtl of control is

begin



    

end architecture;
