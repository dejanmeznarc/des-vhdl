library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use work.screen_pkg.all;

entity sint24 is
  port (
    clk           : in    std_logic;                               -- sistemska ura	
    pin_io_data   : inout std_logic_vector(7 downto 0);            -- IO modul
    pin_io_addr   : out   std_logic_vector(1 downto 0);
    pin_io_clkout : out   std_logic;
    pin_led       : out   unsigned(7 downto 0) := (others => '0'); -- LED
    pin_key       : in    unsigned(1 downto 0)
  );
end entity;

architecture RTL of sint24 is

  signal matrixData     : unsigned(7 downto 0);
  signal buttonData     : unsigned(3 downto 0);
  signal buttonDataPrev : unsigned(3 downto 0);

  signal matrixLine : unsigned(4 downto 0);

  signal counter : unsigned(24 downto 0);
  signal janez   : unsigned(24 downto 0);

  signal offset  : unsigned(2 downto 0) := (others => '0');
  signal offset2 : unsigned(2 downto 0) := (others => '0');

  signal screen : screen_t := (
    "11111",
    "00001",
    "00001",
    "10001",
    "00001",
    "00001",
    "11111"
  );
begin

  identifier: process (clk)
  begin
    if (rising_edge(clk)) then
      counter <= counter + 1;
    end if;
  end process; -- identifier

  interface_inst: entity work.interface
    port map (
      clk      => clk,
      buttons  => buttonData,
      matrix   => matrixData,
      pin_addr => pin_io_addr,
      pin_data => pin_io_data,
      pin_clk  => pin_io_clkout
    );

  matrix_inst: entity work.matrix
    port map (
      clk         => counter(5), -- needs to be at least 4x slower than interface clock
      matrix_data => matrixData,
      screen      => screen
    );

  gpu_driver_inst: entity work.gpu_driver
    port map (
      clk      => counter(24),
      screen   => screen,
      offset_x => offset,
      --offset_y => offset2,
      reset    => not(pin_key(0))
    );

  mikro: process (counter(14), buttonData)
  begin
    if (rising_edge(counter(14))) then

      if (buttonData(0) = '1' and buttonDataPrev(0) = '0') then
        if (offset = 4) then
          offset <= "100";
        else
          offset <= offset + 1;
        end if;
      end if;

      if (buttonData(1) = '1' and buttonDataPrev(1) = '0') then
        if (offset = 0)  then
          offset <= "000";
        else
          offset <= offset - 1;
        end if;
      end if;

      buttonDataPrev <= buttonData;

    end if;



    -- if (not(pin_key(0)) = '1') then
      -- offset <= "010";
    -- end if;
  end process; -- mikro

  pin_led(2 downto 0) <= offset(2 downto 0);

  pin_led(7 downto 5) <= offset2(2 downto 0);

end architecture;
